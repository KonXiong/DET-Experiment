module clock
input 