module Number_Clock;
endmodule